--Universidade Federal de Pelotas--
--Unidade: CDTEC
--Curso: Ciência da computação
--Disciplina: Sistemas Digitais Avançados
--Prof°: Rafael Iankowski Soares
--Aluno: Maicon de Menezes
--Projeto: Trabalho Prático I
--Módulo: Decodificador de 32 Saídas
--Descrição: O código descreve o circuito de um Decodificador de 32 Saídas usado para selecionar qual registrador
--será utilizado para escrita.
library ieee;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
 
entity registerSelector32b is port(
	selectRegister :IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
	registerEnabled:OUT STD_LOGIC_VECTOR (31 DOWNTO 0));
END registerSelector32b;
	
ARCHITECTURE archRegisterSelector32b OF registerSelector32b IS
BEGIN
	WITH selectRegister SELECT
		registerEnabled <= 
		"10000000000000000000000000000000" WHEN "00000",
		"01000000000000000000000000000000" WHEN "00001",
		"00100000000000000000000000000000" WHEN "00010",
		"00010000000000000000000000000000" WHEN "00011",
		"00001000000000000000000000000000" WHEN "00100",
		"00000100000000000000000000000000" WHEN "00101",
		"00000010000000000000000000000000" WHEN "00110",
		"00000001000000000000000000000000" WHEN "00111",
		"00000000100000000000000000000000" WHEN "01000",
		"00000000010000000000000000000000" WHEN "01001",
		"00000000001000000000000000000000" WHEN "01010",
		"00000000000100000000000000000000" WHEN "01011",
		"00000000000010000000000000000000" WHEN "01100",
		"00000000000001000000000000000000" WHEN "01101",
		"00000000000000100000000000000000" WHEN "01110",
		"00000000000000010000000000000000" WHEN "01111",
		"00000000000000001000000000000000" WHEN "10000",
		"00000000000000000100000000000000" WHEN "10001",
		"00000000000000000010000000000000" WHEN "10010",
		"00000000000000000001000000000000" WHEN "10011",
		"00000000000000000000100000000000" WHEN "10100",
		"00000000000000000000010000000000" WHEN "10101",
		"00000000000000000000001000000000" WHEN "10110",
		"00000000000000000000000100000000" WHEN "10111",
		"00000000000000000000000010000000" WHEN "11000",
		"00000000000000000000000001000000" WHEN "11001",
		"00000000000000000000000000100000" WHEN "11010",
		"00000000000000000000000000010000" WHEN "11011",
		"00000000000000000000000000001000" WHEN "11100",
		"00000000000000000000000000000100" WHEN "11101",
		"00000000000000000000000000000010" WHEN "11110",
		"00000000000000000000000000000001" WHEN "11111",
		"00000000000000000000000000000000" WHEN OTHERS;
	END archRegisterSelector32b;